// soon to come, will work for the Intel 3168ngw 
